* SPICE NETLIST
***************************************

.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_vtg_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=2
M0 5 1 3 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=2.282e-13 AS=1.834e-13 PD=3.54e-06 PS=3.49e-06 $X=0 $Y=0 $D=5
M1 4 2 5 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=1.77425e-13 AS=2.282e-13 PD=3.485e-06 PS=3.54e-06 $X=380 $Y=0 $D=5
.ENDS
***************************************
.SUBCKT pmos_vtg_0 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 3 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=2.016e-13 AS=1.512e-13 PD=3.16e-06 PS=3.11e-06 $X=0 $Y=0 $D=4
M1 3 2 4 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=1.58175e-13 AS=2.016e-13 PD=3.105e-06 PS=3.16e-06 $X=380 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT M1_POLY_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X0 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X1 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT M1_N_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_P_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT INVERTER 1 2 3 4
** N=4 EP=4 IP=16 FDC=2
M0 3 4 1 1 NMOS_VTG L=5e-08 W=1.44e-06 AD=1.161e-13 AS=1.0845e-13 PD=3.36e-06 PS=3.19e-06 $X=2045 $Y=110 $D=5
M1 3 4 2 2 PMOS_VTG L=5e-08 W=1.96e-06 AD=1.6015e-13 AS=1.57e-13 PD=4.57e-06 PS=4.5e-06 $X=2040 $Y=3340 $D=4
.ENDS
***************************************
.SUBCKT MUX 1 2 3 4 5 6
** N=9 EP=6 IP=19 FDC=14
X0 4 1 3 7 9 NAND $T=3445 -2060 0 0 $X=3990 $Y=2225
X1 9 1 3 5 2 NAND $T=4660 -2060 0 0 $X=5205 $Y=2225
X2 7 1 3 6 8 NAND $T=5875 -2060 0 0 $X=6420 $Y=2225
X3 1 3 8 2 INVERTER $T=6025 2225 0 0 $X=7635 $Y=2225
.ENDS
***************************************
.SUBCKT NAND_0 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X0 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X1 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT XOR 1 2 3 4 5
** N=9 EP=5 IP=23 FDC=16
X0 2 4 6 1 INVERTER $T=2780 740 1 180 $X=295 $Y=740
X1 2 4 8 3 INVERTER $T=3335 740 0 0 $X=4945 $Y=740
X2 7 2 4 3 6 NAND_0 $T=755 -3545 0 0 $X=1300 $Y=740
X3 5 2 4 7 9 NAND_0 $T=1970 -3545 0 0 $X=2515 $Y=740
X4 9 2 4 1 8 NAND_0 $T=3185 -3545 0 0 $X=3730 $Y=740
.ENDS
***************************************
.SUBCKT NOR 1 2 3 4 5
** N=6 EP=5 IP=4 FDC=4
M0 1 4 3 1 NMOS_VTG L=5e-08 W=7.2e-07 AD=1.008e-13 AS=5.85e-14 PD=1.72e-06 PS=1.76e-06 $X=3705 $Y=545 $D=5
M1 3 5 1 1 NMOS_VTG L=5e-08 W=7.2e-07 AD=5.31e-14 AS=1.008e-13 PD=1.64e-06 PS=1.72e-06 $X=4085 $Y=545 $D=5
M2 6 4 2 2 PMOS_VTG L=5e-08 W=1.56e-06 AD=2.184e-13 AS=1.515e-13 PD=3.4e-06 PS=3.32e-06 $X=3705 $Y=2345 $D=4
M3 3 5 6 2 PMOS_VTG L=5e-08 W=1.56e-06 AD=1.4625e-13 AS=2.184e-13 PD=3.32e-06 PS=3.4e-06 $X=4085 $Y=2345 $D=4
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=8
X0 2 4 5 1 3 NAND_0 $T=0 0 0 0 $X=545 $Y=4285
X1 7 4 5 6 8 NAND_0 $T=1215 0 0 0 $X=1760 $Y=4285
.ENDS
***************************************
.SUBCKT M3_M2_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFF 1 2 3 4 5 6
** N=12 EP=6 IP=42 FDC=30
X8 1 3 11 12 INVERTER $T=1475 1060 0 0 $X=3085 $Y=1060
X9 12 1 3 10 8 NAND_0 $T=3500 -3225 1 180 $X=1740 $Y=1060
X10 10 7 8 1 3 9 8 6 ICV_2 $T=-6095 -3225 0 0 $X=-5550 $Y=1060
X11 10 2 4 1 3 2 4 9 ICV_2 $T=-3665 -3225 0 0 $X=-3120 $Y=1060
X12 7 10 5 1 3 5 9 11 ICV_2 $T=-1235 -3225 0 0 $X=-690 $Y=1060
.ENDS
***************************************
.SUBCKT FA 1 2 3 4 5 6 7
** N=10 EP=7 IP=25 FDC=44
X0 8 3 5 1 2 NAND_0 $T=9190 -2010 0 0 $X=9735 $Y=2275
X1 6 3 5 8 10 NAND_0 $T=10405 -2010 0 0 $X=10950 $Y=2275
X2 10 3 5 4 9 NAND_0 $T=11620 -2010 0 0 $X=12165 $Y=2275
X3 2 3 1 5 9 XOR $T=13080 1535 0 0 $X=13375 $Y=2275
X4 4 3 9 5 7 XOR $T=18760 1535 0 0 $X=19055 $Y=2275
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=60
X0 8 3 1 4 9 2 DFF $T=0 0 0 0 $X=-5550 $Y=1060
X1 8 6 1 7 9 5 DFF $T=9640 0 0 0 $X=4090 $Y=1060
.ENDS
***************************************
.SUBCKT ICV_4
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=12 FDC=28
X0 2 9 5 1 3 4 MUX $T=0 0 0 0 $X=3990 $Y=2225
X1 2 10 5 6 7 8 MUX $T=4650 0 0 0 $X=8640 $Y=2225
.ENDS
***************************************
.SUBCKT MULT 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
** N=25 EP=15 IP=89 FDC=176
X8 4 7 6 17 3 4 MUX $T=6560 -1025 0 0 $X=10550 $Y=1200
X9 4 7 6 25 4 5 MUX $T=50840 -1025 0 0 $X=54830 $Y=1200
X10 18 4 6 7 8 NAND_0 $T=14655 -3085 0 0 $X=15200 $Y=1200
X11 23 4 6 8 9 NAND_0 $T=43770 -3085 0 0 $X=44315 $Y=1200
X17 10 4 17 16 6 16 1 2 18 14 ICV_5 $T=-2740 -1025 0 0 $X=1250 $Y=1200
X18 11 4 20 19 6 19 4 3 15 18 ICV_5 $T=12425 -1025 0 0 $X=16415 $Y=1200
X19 20 4 1 5 6 12 22 21 7 15 ICV_5 $T=21725 -1025 0 0 $X=25715 $Y=1200
X20 21 4 4 5 6 22 3 2 23 7 ICV_5 $T=31025 -1025 0 0 $X=35015 $Y=1200
X21 13 4 25 24 6 24 2 1 23 14 ICV_5 $T=41540 -1025 0 0 $X=45530 $Y=1200
.ENDS
***************************************
.SUBCKT CALC vdd! gnd! I0 I1 I2 I3 B00 B10 B20 B30 S00 S10 O0 O1 O2 O3 S2 CLK
** N=64 EP=18 IP=234 FDC=832
X27 gnd! vdd! 47 46 INVERTER $T=88195 2275 0 0 $X=89805 $Y=2275
X28 gnd! S2 vdd! 4 I0 3 MUX $T=-19560 -7785 1 180 $X=-28075 $Y=-5560
X29 gnd! S2 vdd! 7 I1 6 MUX $T=-5270 -7785 1 180 $X=-13785 $Y=-5560
X30 gnd! S2 vdd! 10 I2 9 MUX $T=9020 -7785 1 180 $X=505 $Y=-5560
X31 gnd! S2 vdd! 13 I3 12 MUX $T=23310 -7785 1 180 $X=14795 $Y=-5560
X32 gnd! 28 vdd! 53 52 24 MUX $T=37515 50 0 0 $X=41505 $Y=2275
X33 gnd! 28 vdd! 27 26 18 MUX $T=65015 50 0 0 $X=69005 $Y=2275
X34 gnd! 59 vdd! 3 2 14 MUX $T=91015 -7785 0 0 $X=95005 $Y=-5560
X35 gnd! 28 vdd! 56 32 21 MUX $T=93650 50 0 0 $X=97640 $Y=2275
X36 gnd! 59 vdd! 6 5 20 MUX $T=95665 -7785 0 0 $X=99655 $Y=-5560
X37 gnd! 59 vdd! 9 8 30 MUX $T=100315 -7785 0 0 $X=104305 $Y=-5560
X38 gnd! 59 vdd! 12 31 34 MUX $T=104965 -7785 0 0 $X=108955 $Y=-5560
X39 23 gnd! O0 vdd! 14 XOR $T=29885 1535 0 0 $X=30180 $Y=2275
X40 23 gnd! 24 vdd! 52 XOR $T=35555 1535 0 0 $X=35850 $Y=2275
X41 25 gnd! 19 vdd! 26 XOR $T=63055 1535 0 0 $X=63350 $Y=2275
X42 55 gnd! 22 vdd! 32 XOR $T=91690 1535 0 0 $X=91985 $Y=2275
X43 56 gnd! O3 vdd! 33 XOR $T=102010 1535 0 0 $X=102305 $Y=2275
X44 33 gnd! 29 vdd! 34 XOR $T=107675 1535 0 0 $X=107970 $Y=2275
X45 gnd! vdd! 54 15 16 NOR $T=42685 1840 0 0 $X=46080 $Y=2275
X46 gnd! vdd! 25 23 24 NOR $T=58705 1840 0 0 $X=62100 $Y=2275
X47 gnd! vdd! 46 23 24 NOR $T=85160 1840 0 0 $X=88555 $Y=2275
X48 gnd! vdd! 55 47 18 NOR $T=87340 1840 0 0 $X=90735 $Y=2275
X56 gnd! O0 vdd! 15 CLK 4 DFF $T=-17870 -6620 0 0 $X=-23420 $Y=-5560
X57 gnd! O1 vdd! 57 CLK 7 DFF $T=-3580 -6620 0 0 $X=-9130 $Y=-5560
X58 gnd! O2 vdd! 58 CLK 10 DFF $T=10710 -6620 0 0 $X=5160 $Y=-5560
X59 gnd! 59 vdd! 60 CLK S10 DFF $T=82840 -6620 0 0 $X=77290 $Y=-5560
X60 53 O1 gnd! 54 vdd! 17 20 FA $T=37465 0 0 0 $X=47200 $Y=2275
X61 27 O2 gnd! 17 vdd! 29 30 FA $T=63920 0 0 0 $X=73655 $Y=2275
X62 vdd! 13 O3 61 B00 23 16 gnd! CLK ICV_3 $T=25000 -6620 0 0 $X=19450 $Y=-5560
X63 vdd! B10 24 62 B20 18 19 gnd! CLK ICV_3 $T=44280 -6620 0 0 $X=38730 $Y=-5560
X64 vdd! B30 21 22 S00 28 11 gnd! CLK ICV_3 $T=63560 -6620 0 0 $X=58010 $Y=-5560
X65 O2 O1 O3 gnd! O0 vdd! 28 22 11 2 5 8 31 18 24 MULT $T=-29315 1075 0 0 $X=-28065 $Y=2275
.ENDS
***************************************
