* SPICE NETLIST
***************************************

.SUBCKT M1_POLY_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_N_3
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_P_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT Inverter gnd! vdd! Out In
** N=4 EP=4 IP=16 FDC=2
M0 Out In gnd! gnd! NMOS_VTG L=5e-08 W=1.44e-06 AD=1.161e-13 AS=1.0845e-13 PD=3.36e-06 PS=3.19e-06 $X=2045 $Y=110 $D=5
M1 Out In vdd! vdd! PMOS_VTG L=5e-08 W=1.96e-06 AD=1.6015e-13 AS=1.57e-13 PD=4.57e-06 PS=4.5e-06 $X=2040 $Y=3340 $D=4
.ENDS
***************************************
.SUBCKT OR gnd! vdd! 3 A B Output
** N=7 EP=6 IP=8 FDC=6
M0 gnd! A 3 gnd! NMOS_VTG L=5e-08 W=7.2e-07 AD=1.008e-13 AS=5.85e-14 PD=1.72e-06 PS=1.76e-06 $X=-815 $Y=-1620 $D=5
M1 3 B gnd! gnd! NMOS_VTG L=5e-08 W=7.2e-07 AD=5.31e-14 AS=1.008e-13 PD=1.64e-06 PS=1.72e-06 $X=-435 $Y=-1620 $D=5
M2 7 A vdd! vdd! PMOS_VTG L=5e-08 W=1.56e-06 AD=2.184e-13 AS=1.515e-13 PD=3.4e-06 PS=3.32e-06 $X=-815 $Y=180 $D=4
M3 3 B 7 vdd! PMOS_VTG L=5e-08 W=1.56e-06 AD=1.4625e-13 AS=2.184e-13 PD=3.32e-06 PS=3.4e-06 $X=-435 $Y=180 $D=4
X8 gnd! vdd! Output 3 Inverter $T=-1475 -3170 0 0 $X=135 $Y=-3170
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9
** N=10 EP=9 IP=12 FDC=12
X0 4 5 3 1 2 6 OR $T=0 0 0 0 $X=-1125 $Y=-3170
X1 4 5 10 7 8 9 OR $T=2190 0 0 0 $X=1065 $Y=-3170
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
** N=16 EP=15 IP=18 FDC=24
X0 1 2 16 3 4 5 6 7 8 ICV_2 $T=0 0 0 0 $X=-1125 $Y=-3170
X1 9 10 11 3 4 12 13 14 15 ICV_2 $T=0 7820 0 0 $X=-1125 $Y=4650
.ENDS
***************************************
.SUBCKT dcont_8
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_vtg_0 1 2 3 4
** N=4 EP=4 IP=2 FDC=1
M0 2 3 1 4 NMOS_VTG L=5e-08 W=2.8e-07 AD=2.94e-14 AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 $X=0 $Y=0 $D=5
.ENDS
***************************************
.SUBCKT pmos_vtg_1 1 2 3 4
** N=4 EP=4 IP=2 FDC=1
M0 2 3 1 4 PMOS_VTG L=5e-08 W=3e-07 AD=3.15e-14 AS=3.15e-14 PD=8.1e-07 PS=8.1e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT XOR B Output A 4 5 6 7
** N=8 EP=7 IP=28 FDC=6
X4 4 8 A 6 nmos_vtg_0 $T=2400 2225 0 0 $X=2080 $Y=2115
X5 8 Output B 6 nmos_vtg_0 $T=3140 2225 0 0 $X=2820 $Y=2115
X6 Output B 8 6 nmos_vtg_0 $T=3880 2225 0 0 $X=3560 $Y=2115
X7 5 8 A 7 pmos_vtg_1 $T=2400 3215 0 0 $X=2080 $Y=3105
X8 A Output B 7 pmos_vtg_1 $T=3140 3215 0 0 $X=2820 $Y=3105
X9 Output B A 7 pmos_vtg_1 $T=3880 3215 0 0 $X=3560 $Y=3105
.ENDS
***************************************
.SUBCKT FULL_ADDER_noCOUT gnd! vdd! B A Cin S 7 8
** N=9 EP=8 IP=14 FDC=12
X0 B 9 A gnd! vdd! 7 8 XOR $T=2040 540 0 0 $X=4120 $Y=2435
X1 Cin S 9 gnd! vdd! 7 8 XOR $T=10640 540 1 180 $X=6340 $Y=2435
.ENDS
***************************************
.SUBCKT AND gnd! vdd! B A Output
** N=7 EP=5 IP=6 FDC=6
M0 7 B gnd! gnd! NMOS_VTG L=5e-08 W=1.63e-06 AD=2.282e-13 AS=1.77425e-13 PD=3.54e-06 PS=3.485e-06 $X=-1025 $Y=-3500 $D=5
M1 6 A 7 gnd! NMOS_VTG L=5e-08 W=1.63e-06 AD=1.834e-13 AS=2.282e-13 PD=3.49e-06 PS=3.54e-06 $X=-645 $Y=-3500 $D=5
M2 6 B vdd! vdd! PMOS_VTG L=5e-08 W=1.44e-06 AD=2.016e-13 AS=1.58175e-13 PD=3.16e-06 PS=3.105e-06 $X=-1025 $Y=150 $D=4
M3 vdd! A 6 vdd! PMOS_VTG L=5e-08 W=1.44e-06 AD=1.512e-13 AS=2.016e-13 PD=3.11e-06 PS=3.16e-06 $X=-645 $Y=150 $D=4
X6 gnd! vdd! Output 6 Inverter $T=-1610 -4155 0 0 $X=0 $Y=-4155
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=12
X0 1 2 3 4 5 AND $T=0 0 0 0 $X=-1360 $Y=-4155
X1 1 2 6 7 8 AND $T=2230 0 0 0 $X=870 $Y=-4155
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=16 FDC=24
X0 1 2 3 4 5 6 7 8 ICV_4 $T=0 0 0 0 $X=-1360 $Y=-4155
X1 1 2 9 10 11 12 13 14 ICV_4 $T=0 7820 0 0 $X=-1360 $Y=3665
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26
** N=26 EP=26 IP=28 FDC=48
X0 1 2 3 5 7 9 11 13 4 6 8 10 12 14 ICV_5 $T=0 0 0 0 $X=-1360 $Y=-4155
X1 1 2 15 17 19 21 23 25 16 18 20 22 24 26 ICV_5 $T=4460 0 0 0 $X=3100 $Y=-4155
.ENDS
***************************************
.SUBCKT LOOKAHEAD B<0> A<0> B<1> A<1> B<2> B<6> A<2> A<6> B<3> A<3> B<4> A<4> A<7> B<5> A<5> gnd! vdd! S<0> Cout S<1>
+ S<2> S<3> S<4> S<5> S<6> S<7>
** N=114 EP=26 IP=337 FDC=516
X4 gnd! vdd! 94 11 87 61 OR $T=77350 7335 0 0 $X=76225 $Y=4165
X5 52 88 95 gnd! vdd! 89 50 89 Cout ICV_2 $T=77350 15155 0 0 $X=76225 $Y=11985
X6 A<1> B<1> gnd! vdd! 13 10 14 63 6 61 97 62 27 62 64 ICV_3 $T=42310 7335 0 0 $X=41185 $Y=4165
X7 A<2> B<2> gnd! vdd! 66 39 28 67 22 64 65 98 A<6> B<6> 24 ICV_3 $T=46690 7335 0 0 $X=45565 $Y=4165
X8 25 67 gnd! vdd! 68 A<3> B<3> 34 21 42 99 69 38 69 70 ICV_3 $T=51070 7335 0 0 $X=49945 $Y=4165
X9 32 41 gnd! vdd! 71 37 71 73 36 70 100 72 33 72 74 ICV_3 $T=55450 7335 0 0 $X=54325 $Y=4165
X10 35 73 gnd! vdd! 75 A<4> B<4> 47 29 74 101 76 26 76 77 ICV_3 $T=59830 7335 0 0 $X=58705 $Y=4165
X11 12 8 gnd! vdd! 78 2 78 79 A<7> B<4> 102 48 46 60 80 ICV_3 $T=64210 7335 0 0 $X=63085 $Y=4165
X12 51 79 gnd! vdd! 104 49 82 83 59 80 103 81 58 81 84 ICV_3 $T=68590 7335 0 0 $X=67465 $Y=4165
X13 A<5> 85 gnd! vdd! 4 40 15 87 55 84 105 86 54 86 88 ICV_3 $T=72970 7335 0 0 $X=71845 $Y=4165
X14 gnd! 92 A<0> 113 nmos_vtg_0 $T=23430 1605 0 0 $X=23110 $Y=1495
X15 92 S<0> B<0> 113 nmos_vtg_0 $T=24170 1605 0 0 $X=23850 $Y=1495
X16 S<0> B<0> 92 113 nmos_vtg_0 $T=24910 1605 0 0 $X=24590 $Y=1495
X17 vdd! 92 A<0> 114 pmos_vtg_1 $T=23430 2595 0 0 $X=23110 $Y=2485
X18 A<0> S<0> B<0> 114 pmos_vtg_1 $T=24170 2595 0 0 $X=23850 $Y=2485
X19 S<0> B<0> A<0> 114 pmos_vtg_1 $T=24910 2595 0 0 $X=24590 $Y=2485
X20 gnd! vdd! B<1> A<1> 5 S<1> 113 114 FULL_ADDER_noCOUT $T=21210 -1160 0 0 $X=25330 $Y=1025
X21 gnd! vdd! B<2> A<2> 63 S<2> 113 114 FULL_ADDER_noCOUT $T=25690 -1160 0 0 $X=29810 $Y=1025
X22 gnd! vdd! B<3> A<3> 68 S<3> 113 114 FULL_ADDER_noCOUT $T=30170 -1160 0 0 $X=34290 $Y=1025
X23 gnd! vdd! B<4> A<4> 75 S<4> 113 114 FULL_ADDER_noCOUT $T=34650 -1160 0 0 $X=38770 $Y=1025
X24 gnd! vdd! B<5> A<5> 83 S<5> 113 114 FULL_ADDER_noCOUT $T=39130 -1160 0 0 $X=43250 $Y=1025
X25 gnd! vdd! B<6> A<6> 65 S<6> 113 114 FULL_ADDER_noCOUT $T=43610 -1160 0 0 $X=47730 $Y=1025
X26 gnd! vdd! B<4> A<7> 77 S<7> 113 114 FULL_ADDER_noCOUT $T=48090 -1160 0 0 $X=52210 $Y=1025
X27 gnd! vdd! 49 4 22 51 4 27 42 48 59 21 48 60 ICV_5 $T=38025 8320 0 0 $X=36665 $Y=4165
X28 gnd! vdd! B<0> 2 A<0> 4 5 6 B<1> 8 A<1> 4 10 11 5 12 13 4 14 15
+ B<2> B<6> A<2> A<6> 20 21
+ ICV_6 $T=2345 8320 0 0 $X=985 $Y=4165
X29 gnd! vdd! 14 22 23 24 25 26 10 27 23 24 28 29 B<3> 6 A<3> 24 32 33
+ 25 11 34 24 35 36
+ ICV_6 $T=11265 8320 0 0 $X=9905 $Y=4165
X30 gnd! vdd! 28 15 34 24 37 38 39 40 34 24 41 42 B<4> B<4> A<4> A<7> 12 46
+ 35 26 47 48 49 50
+ ICV_6 $T=20185 8320 0 0 $X=18825 $Y=4165
X31 gnd! vdd! 37 29 47 48 51 52 41 33 47 53 2 54 32 36 47 48 8 55
+ B<5> 38 A<5> 48 40 58
+ ICV_6 $T=29105 8320 0 0 $X=27745 $Y=4165
.ENDS
***************************************
