* SPICE NETLIST
***************************************

.SUBCKT M1_POLY_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_N_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_P_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT INVERTER 1 2 3 4
** N=4 EP=4 IP=16 FDC=2
M0 3 4 1 1 NMOS_VTG L=5e-08 W=1.44e-06 AD=1.161e-13 AS=1.0845e-13 PD=3.36e-06 PS=3.19e-06 $X=2045 $Y=110 $D=5
M1 3 4 2 2 PMOS_VTG L=5e-08 W=1.96e-06 AD=1.6015e-13 AS=1.57e-13 PD=4.57e-06 PS=4.5e-06 $X=2040 $Y=3340 $D=4
.ENDS
***************************************
.SUBCKT nmos_vtg_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=2
M0 5 1 3 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=2.282e-13 AS=1.834e-13 PD=3.54e-06 PS=3.49e-06 $X=0 $Y=0 $D=5
M1 4 2 5 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=1.77425e-13 AS=2.282e-13 PD=3.485e-06 PS=3.54e-06 $X=380 $Y=0 $D=5
.ENDS
***************************************
.SUBCKT pmos_vtg_0 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 3 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=2.016e-13 AS=1.512e-13 PD=3.16e-06 PS=3.11e-06 $X=0 $Y=0 $D=4
M1 3 2 4 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=1.58175e-13 AS=2.016e-13 PD=3.105e-06 PS=3.16e-06 $X=380 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT NAND 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT XOR 2 3 5 7 9
** N=9 EP=5 IP=23 FDC=16
X0 3 7 1 2 INVERTER $T=2780 740 1 180 $X=295 $Y=740
X1 3 7 6 5 INVERTER $T=3335 740 0 0 $X=4945 $Y=740
X2 4 3 7 5 1 NAND $T=755 -3545 0 0 $X=1300 $Y=740
X3 9 3 7 4 8 NAND $T=1970 -3545 0 0 $X=2515 $Y=740
X4 8 3 7 2 6 NAND $T=3185 -3545 0 0 $X=3730 $Y=740
.ENDS
***************************************
.SUBCKT NAND_0 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT ADD2 gnd! S0 A2 C1 B0 B1 vdd! B2 C2 X2 B2N
** N=21 EP=11 IP=53 FDC=78
M0 gnd! B0 1 gnd! NMOS_VTG L=5e-08 W=7.2e-07 AD=1.008e-13 AS=5.85e-14 PD=1.72e-06 PS=1.76e-06 $X=9450 $Y=1770 $D=5
M1 1 B1 gnd! gnd! NMOS_VTG L=5e-08 W=7.2e-07 AD=5.31e-14 AS=1.008e-13 PD=1.64e-06 PS=1.72e-06 $X=9830 $Y=1770 $D=5
M2 21 B0 vdd! vdd! PMOS_VTG L=5e-08 W=1.56e-06 AD=2.184e-13 AS=1.515e-13 PD=3.4e-06 PS=3.32e-06 $X=9450 $Y=3570 $D=4
M3 1 B1 21 vdd! PMOS_VTG L=5e-08 W=1.56e-06 AD=1.4625e-13 AS=2.184e-13 PD=3.32e-06 PS=3.4e-06 $X=9830 $Y=3570 $D=4
X8 gnd! vdd! 7 S0 INVERTER $T=18080 1660 0 0 $X=19690 $Y=1660
X9 8 gnd! vdd! 3 A2 NAND $T=20150 -2625 0 0 $X=20695 $Y=1660
X10 C2 gnd! vdd! 8 18 NAND $T=21365 -2625 0 0 $X=21910 $Y=1660
X11 18 gnd! vdd! C1 11 NAND $T=22580 -2625 0 0 $X=23125 $Y=1660
X12 1 gnd! B2N vdd! 2 XOR $T=10095 920 0 0 $X=10390 $Y=1660
X13 A2 gnd! 3 vdd! 11 XOR $T=24040 920 0 0 $X=24335 $Y=1660
X14 C1 gnd! 11 vdd! X2 XOR $T=29720 920 0 0 $X=30015 $Y=1660
X15 3 gnd! vdd! 4 15 NAND_0 $T=15500 -2625 0 0 $X=16045 $Y=1660
X16 15 gnd! vdd! 2 S0 NAND_0 $T=16715 -2625 0 0 $X=17260 $Y=1660
X17 4 gnd! vdd! B2 7 NAND_0 $T=17930 -2625 0 0 $X=18475 $Y=1660
.ENDS
***************************************
