* SPICE NETLIST
***************************************

.SUBCKT M1_N_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_P_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT M1_POLY_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVERTER 1 2 3 4
** N=4 EP=4 IP=16 FDC=2
M0 3 4 1 1 NMOS_VTG L=5e-08 W=1.44e-06 AD=1.161e-13 AS=1.0845e-13 PD=3.36e-06 PS=3.19e-06 $X=2045 $Y=110 $D=5
M1 3 4 2 2 PMOS_VTG L=5e-08 W=1.96e-06 AD=1.6015e-13 AS=1.57e-13 PD=4.57e-06 PS=4.5e-06 $X=2040 $Y=3340 $D=4
.ENDS
***************************************
.SUBCKT nmos_vtg_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=2
M0 5 1 3 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=2.282e-13 AS=1.834e-13 PD=3.54e-06 PS=3.49e-06 $X=0 $Y=0 $D=5
M1 4 2 5 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=1.77425e-13 AS=2.282e-13 PD=3.485e-06 PS=3.54e-06 $X=380 $Y=0 $D=5
.ENDS
***************************************
.SUBCKT pmos_vtg_0 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 3 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=2.016e-13 AS=1.512e-13 PD=3.16e-06 PS=3.11e-06 $X=0 $Y=0 $D=4
M1 3 2 4 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=1.58175e-13 AS=2.016e-13 PD=3.105e-06 PS=3.16e-06 $X=380 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT NAND 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT XOR 1 2 3 4 5
** N=9 EP=5 IP=23 FDC=16
X0 2 4 6 1 INVERTER $T=2780 740 1 180 $X=295 $Y=740
X1 2 4 8 3 INVERTER $T=3335 740 0 0 $X=4945 $Y=740
X2 7 2 4 3 6 NAND $T=755 -3545 0 0 $X=1300 $Y=740
X3 5 2 4 7 9 NAND $T=1970 -3545 0 0 $X=2515 $Y=740
X4 9 2 4 1 8 NAND $T=3185 -3545 0 0 $X=3730 $Y=740
.ENDS
***************************************
.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND_0 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT ADD1
** N=20 EP=0 IP=59 FDC=78
M0 2 13 8 2 NMOS_VTG L=5e-08 W=7.2e-07 AD=1.008e-13 AS=5.85e-14 PD=1.72e-06 PS=1.76e-06 $X=40000 $Y=-10795 $D=5
M1 8 14 2 2 NMOS_VTG L=5e-08 W=7.2e-07 AD=5.31e-14 AS=1.008e-13 PD=1.64e-06 PS=1.72e-06 $X=40380 $Y=-10795 $D=5
M2 20 13 10 10 PMOS_VTG L=5e-08 W=1.56e-06 AD=2.184e-13 AS=1.515e-13 PD=3.4e-06 PS=3.32e-06 $X=40000 $Y=-8995 $D=4
M3 8 14 20 10 PMOS_VTG L=5e-08 W=1.56e-06 AD=1.4625e-13 AS=2.184e-13 PD=3.32e-06 PS=3.4e-06 $X=40380 $Y=-8995 $D=4
X8 2 10 4 3 INVERTER $T=37150 -10905 0 0 $X=38760 $Y=-10905
X9 5 2 10 6 7 NAND $T=40265 -15190 0 0 $X=40810 $Y=-10905
X10 15 2 10 5 12 NAND $T=41480 -15190 0 0 $X=42025 $Y=-10905
X11 12 2 10 8 9 NAND $T=42695 -15190 0 0 $X=43240 $Y=-10905
X12 19 2 18 10 16 XOR $T=29165 -11645 0 0 $X=29460 $Y=-10905
X13 7 2 6 10 9 XOR $T=44155 -11645 0 0 $X=44450 $Y=-10905
X14 8 2 9 10 17 XOR $T=49835 -11645 0 0 $X=50130 $Y=-10905
X21 6 2 10 1 11 NAND_0 $T=34570 -15190 0 0 $X=35115 $Y=-10905
X22 11 2 10 16 3 NAND_0 $T=35785 -15190 0 0 $X=36330 $Y=-10905
X23 1 2 10 18 4 NAND_0 $T=37000 -15190 0 0 $X=37545 $Y=-10905
.ENDS
***************************************
