* SPICE NETLIST
***************************************

.SUBCKT M1_POLY_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_N_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR 1 2 3 4
** N=6 EP=4 IP=4 FDC=4
M0 1 4 3 1 NMOS_VTG L=5e-08 W=7.2e-07 AD=1.008e-13 AS=5.85e-14 PD=1.72e-06 PS=1.76e-06 $X=3705 $Y=545 $D=5
M1 3 5 1 1 NMOS_VTG L=5e-08 W=7.2e-07 AD=5.31e-14 AS=1.008e-13 PD=1.64e-06 PS=1.72e-06 $X=4085 $Y=545 $D=5
M2 6 4 2 2 PMOS_VTG L=5e-08 W=1.56e-06 AD=2.184e-13 AS=1.515e-13 PD=3.4e-06 PS=3.32e-06 $X=3705 $Y=2345 $D=4
M3 3 5 6 2 PMOS_VTG L=5e-08 W=1.56e-06 AD=1.4625e-13 AS=2.184e-13 PD=3.32e-06 PS=3.4e-06 $X=4085 $Y=2345 $D=4
.ENDS
***************************************
.SUBCKT M1_P_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT INVERTER 1 2 3 4
** N=4 EP=4 IP=16 FDC=2
M0 3 4 1 1 NMOS_VTG L=5e-08 W=1.44e-06 AD=1.161e-13 AS=1.0845e-13 PD=3.36e-06 PS=3.19e-06 $X=2045 $Y=110 $D=5
M1 3 4 2 2 PMOS_VTG L=5e-08 W=1.96e-06 AD=1.6015e-13 AS=1.57e-13 PD=4.57e-06 PS=4.5e-06 $X=2040 $Y=3340 $D=4
.ENDS
***************************************
.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_vtg_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=2
M0 5 1 3 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=2.282e-13 AS=1.834e-13 PD=3.54e-06 PS=3.49e-06 $X=0 $Y=0 $D=5
M1 4 2 5 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=1.77425e-13 AS=2.282e-13 PD=3.485e-06 PS=3.54e-06 $X=380 $Y=0 $D=5
.ENDS
***************************************
.SUBCKT pmos_vtg_0 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 3 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=2.016e-13 AS=1.512e-13 PD=3.16e-06 PS=3.11e-06 $X=0 $Y=0 $D=4
M1 3 2 4 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=1.58175e-13 AS=2.016e-13 PD=3.105e-06 PS=3.16e-06 $X=380 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT NAND 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT XOR 1 2 3 4
** N=9 EP=4 IP=23 FDC=16
X0 2 3 5 1 INVERTER $T=2780 740 1 180 $X=295 $Y=740
X1 2 3 8 7 INVERTER $T=3335 740 0 0 $X=4945 $Y=740
X2 6 2 3 7 5 NAND $T=755 -3545 0 0 $X=1300 $Y=740
X3 4 2 3 6 9 NAND $T=1970 -3545 0 0 $X=2515 $Y=740
X4 9 2 3 1 8 NAND $T=3185 -3545 0 0 $X=3730 $Y=740
.ENDS
***************************************
.SUBCKT NAND_0 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT ADD3
** N=15 EP=0 IP=46 FDC=72
X0 3 8 7 11 NOR $T=36300 -5670 0 0 $X=39695 $Y=-5235
X1 3 8 12 9 NOR $T=38480 -5670 0 0 $X=41875 $Y=-5235
X2 3 8 9 7 INVERTER $T=39335 -5235 0 0 $X=40945 $Y=-5235
X3 3 8 5 4 INVERTER $T=50815 -5235 0 0 $X=52425 $Y=-5235
X7 12 3 8 1 XOR $T=42830 -5975 0 0 $X=43125 $Y=-5235
X8 13 3 8 6 XOR $T=53150 -5975 0 0 $X=53445 $Y=-5235
X9 6 3 8 14 XOR $T=58815 -5975 0 0 $X=59110 $Y=-5235
X10 13 3 8 2 10 NAND_0 $T=48235 -9520 0 0 $X=48780 $Y=-5235
X11 10 3 8 1 4 NAND_0 $T=49450 -9520 0 0 $X=49995 $Y=-5235
X12 2 3 8 15 5 NAND_0 $T=50665 -9520 0 0 $X=51210 $Y=-5235
.ENDS
***************************************
