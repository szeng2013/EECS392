* SPICE NETLIST
***************************************

.SUBCKT M1_N_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_P_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT M1_POLY_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVERTER 1 2 3 4
** N=4 EP=4 IP=16 FDC=2
M0 3 4 1 1 NMOS_VTG L=5e-08 W=1.44e-06 AD=1.161e-13 AS=1.0845e-13 PD=3.36e-06 PS=3.19e-06 $X=2045 $Y=110 $D=5
M1 3 4 2 2 PMOS_VTG L=5e-08 W=1.96e-06 AD=1.6015e-13 AS=1.57e-13 PD=4.57e-06 PS=4.5e-06 $X=2040 $Y=3340 $D=4
.ENDS
***************************************
.SUBCKT nmos_vtg_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=2
M0 5 1 3 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=2.282e-13 AS=1.834e-13 PD=3.54e-06 PS=3.49e-06 $X=0 $Y=0 $D=5
M1 4 2 5 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=1.77425e-13 AS=2.282e-13 PD=3.485e-06 PS=3.54e-06 $X=380 $Y=0 $D=5
.ENDS
***************************************
.SUBCKT pmos_vtg_0 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 3 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=2.016e-13 AS=1.512e-13 PD=3.16e-06 PS=3.11e-06 $X=0 $Y=0 $D=4
M1 3 2 4 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=1.58175e-13 AS=2.016e-13 PD=3.105e-06 PS=3.16e-06 $X=380 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT NAND 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT XOR 2 3 5 7 9
** N=9 EP=5 IP=23 FDC=16
X0 3 7 1 2 INVERTER $T=2780 740 1 180 $X=295 $Y=740
X1 3 7 6 5 INVERTER $T=3335 740 0 0 $X=4945 $Y=740
X2 4 3 7 5 1 NAND $T=755 -3545 0 0 $X=1300 $Y=740
X3 9 3 7 4 8 NAND $T=1970 -3545 0 0 $X=2515 $Y=740
X4 8 3 7 2 6 NAND $T=3185 -3545 0 0 $X=3730 $Y=740
.ENDS
***************************************
.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND_0 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT MUX 2 3 6 7 8 9
** N=9 EP=6 IP=19 FDC=14
X0 2 6 4 3 INVERTER $T=6025 2225 0 0 $X=7635 $Y=2225
X1 7 2 6 1 5 NAND_0 $T=3445 -2060 0 0 $X=3990 $Y=2225
X2 5 2 6 8 3 NAND_0 $T=4660 -2060 0 0 $X=5205 $Y=2225
X3 1 2 6 9 4 NAND_0 $T=5875 -2060 0 0 $X=6420 $Y=2225
.ENDS
***************************************
.SUBCKT NOR 1 2 3 4 5
** N=6 EP=5 IP=4 FDC=4
M0 1 4 3 1 NMOS_VTG L=5e-08 W=7.2e-07 AD=1.008e-13 AS=5.85e-14 PD=1.72e-06 PS=1.76e-06 $X=3705 $Y=545 $D=5
M1 3 5 1 1 NMOS_VTG L=5e-08 W=7.2e-07 AD=5.31e-14 AS=1.008e-13 PD=1.64e-06 PS=1.72e-06 $X=4085 $Y=545 $D=5
M2 6 4 2 2 PMOS_VTG L=5e-08 W=1.56e-06 AD=2.184e-13 AS=1.515e-13 PD=3.4e-06 PS=3.32e-06 $X=3705 $Y=2345 $D=4
M3 3 5 6 2 PMOS_VTG L=5e-08 W=1.56e-06 AD=1.4625e-13 AS=2.184e-13 PD=3.32e-06 PS=3.4e-06 $X=4085 $Y=2345 $D=4
.ENDS
***************************************
.SUBCKT FA 2 3 4 5 7 9 10
** N=10 EP=7 IP=25 FDC=44
X0 1 4 7 2 3 NAND $T=9190 -2010 0 0 $X=9735 $Y=2275
X1 9 4 7 1 8 NAND $T=10405 -2010 0 0 $X=10950 $Y=2275
X2 8 4 7 5 6 NAND $T=11620 -2010 0 0 $X=12165 $Y=2275
X3 3 4 2 7 6 XOR $T=13080 1535 0 0 $X=13375 $Y=2275
X4 5 4 6 7 10 XOR $T=18760 1535 0 0 $X=19055 $Y=2275
.ENDS
***************************************
.SUBCKT ADDER B0 B1 B2 X0 vdd! A0N B0N X1 gnd! X2 B3 X3 A0 S0 B2N B3N A3 A1 A2
** N=33 EP=19 IP=95 FDC=244
X0 gnd! vdd! 19 18 INVERTER $T=62255 1585 0 0 $X=63865 $Y=1585
X1 B0 gnd! A0 vdd! X0 XOR $T=3945 845 0 0 $X=4240 $Y=1585
X2 B0 gnd! B1 vdd! 22 XOR $T=9615 845 0 0 $X=9910 $Y=1585
X3 4 gnd! B2N vdd! 5 XOR $T=37115 845 0 0 $X=37410 $Y=1585
X4 25 gnd! B3N vdd! 9 XOR $T=65750 845 0 0 $X=66045 $Y=1585
X5 26 gnd! A3 vdd! 10 XOR $T=76070 845 0 0 $X=76365 $Y=1585
X6 10 gnd! 8 vdd! X3 XOR $T=81735 845 0 0 $X=82030 $Y=1585
X16 gnd! S0 vdd! 23 22 B1 MUX $T=11575 -640 0 0 $X=15565 $Y=1585
X17 gnd! S0 vdd! 6 5 B2 MUX $T=39075 -640 0 0 $X=43065 $Y=1585
X18 gnd! S0 vdd! 26 9 B3 MUX $T=67710 -640 0 0 $X=71700 $Y=1585
X19 gnd! vdd! 24 A0N B0N NOR $T=16745 1150 0 0 $X=20140 $Y=1585
X20 gnd! vdd! 4 B0 B1 NOR $T=32765 1150 0 0 $X=36160 $Y=1585
X21 gnd! vdd! 18 B0 B1 NOR $T=59220 1150 0 0 $X=62615 $Y=1585
X22 gnd! vdd! 25 19 B2 NOR $T=61400 1150 0 0 $X=64795 $Y=1585
X23 23 A1 gnd! 24 vdd! 1 X1 FA $T=11525 -690 0 0 $X=21260 $Y=1585
X24 6 A2 gnd! 1 vdd! 8 X2 FA $T=37980 -690 0 0 $X=47715 $Y=1585
.ENDS
***************************************
