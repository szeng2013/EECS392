* SPICE NETLIST
***************************************

.SUBCKT M1_N_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_P_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT M1_POLY_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND 1 2 3 4 5
** N=6 EP=5 IP=2 FDC=4
M0 6 4 1 2 NMOS_VTG L=5e-08 W=1.63e-06 AD=2.282e-13 AS=1.834e-13 PD=3.54e-06 PS=3.49e-06 $X=945 $Y=4395 $D=5
M1 2 5 6 2 NMOS_VTG L=5e-08 W=1.63e-06 AD=1.77425e-13 AS=2.282e-13 PD=3.485e-06 PS=3.54e-06 $X=1325 $Y=4395 $D=5
M2 1 4 3 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=2.016e-13 AS=1.512e-13 PD=3.16e-06 PS=3.11e-06 $X=945 $Y=8045 $D=4
M3 3 5 1 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=1.58175e-13 AS=2.016e-13 PD=3.105e-06 PS=3.16e-06 $X=1325 $Y=8045 $D=4
.ENDS
***************************************
.SUBCKT MUX 2 3 6 7 8 9
** N=9 EP=6 IP=31 FDC=14
M0 4 3 2 2 NMOS_VTG L=5e-08 W=1.44e-06 AD=1.161e-13 AS=1.0845e-13 PD=3.36e-06 PS=3.19e-06 $X=8070 $Y=2335 $D=5
M1 4 3 6 6 PMOS_VTG L=5e-08 W=1.96e-06 AD=1.6015e-13 AS=1.57e-13 PD=4.57e-06 PS=4.5e-06 $X=8065 $Y=5565 $D=4
X18 7 2 6 1 5 NAND $T=3445 -2060 0 0 $X=3990 $Y=2225
X19 5 2 6 8 3 NAND $T=4660 -2060 0 0 $X=5205 $Y=2225
X20 1 2 6 9 4 NAND $T=5875 -2060 0 0 $X=6420 $Y=2225
.ENDS
***************************************
.SUBCKT OUTPUT O0 Y0 X0 O1 vdd! Y1 X1 O2 Y2 X2 O3 Y3 X3 gnd! S1
** N=15 EP=15 IP=24 FDC=56
X0 gnd! S1 vdd! O0 Y0 X0 MUX $T=-1875 -1380 0 0 $X=2115 $Y=845
X1 gnd! S1 vdd! O1 Y1 X1 MUX $T=2775 -1380 0 0 $X=6765 $Y=845
X2 gnd! S1 vdd! O2 Y2 X2 MUX $T=7425 -1380 0 0 $X=11415 $Y=845
X3 gnd! S1 vdd! O3 Y3 X3 MUX $T=12075 -1380 0 0 $X=16065 $Y=845
.ENDS
***************************************
