* SPICE NETLIST
***************************************

.SUBCKT M1_N_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_P_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT M1_POLY_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVERTER 1 2 3 4
** N=4 EP=4 IP=16 FDC=2
M0 3 4 1 1 NMOS_VTG L=5e-08 W=1.44e-06 AD=1.161e-13 AS=1.0845e-13 PD=3.36e-06 PS=3.19e-06 $X=2045 $Y=110 $D=5
M1 3 4 2 2 PMOS_VTG L=5e-08 W=1.96e-06 AD=1.6015e-13 AS=1.57e-13 PD=4.57e-06 PS=4.5e-06 $X=2040 $Y=3340 $D=4
.ENDS
***************************************
.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_vtg_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=2
M0 5 1 3 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=2.282e-13 AS=1.834e-13 PD=3.54e-06 PS=3.49e-06 $X=0 $Y=0 $D=5
M1 4 2 5 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=1.77425e-13 AS=2.282e-13 PD=3.485e-06 PS=3.54e-06 $X=380 $Y=0 $D=5
.ENDS
***************************************
.SUBCKT pmos_vtg_0 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 3 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=2.016e-13 AS=1.512e-13 PD=3.16e-06 PS=3.11e-06 $X=0 $Y=0 $D=4
M1 3 2 4 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=1.58175e-13 AS=2.016e-13 PD=3.105e-06 PS=3.16e-06 $X=380 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT NAND 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=8
X0 1 5 2 3 4 NAND $T=0 0 0 0 $X=545 $Y=4285
X1 6 5 2 7 8 NAND $T=1215 0 0 0 $X=1760 $Y=4285
.ENDS
***************************************
.SUBCKT M3_M2_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFF 1 2 3 4
** N=12 EP=4 IP=42 FDC=30
X0 1 2 10 12 INVERTER $T=1475 1060 0 0 $X=3085 $Y=1060
X9 12 1 2 9 6 NAND $T=3500 -3225 1 180 $X=1740 $Y=1060
X10 5 2 9 6 1 6 7 4 ICV_2 $T=-6095 -3225 0 0 $X=-5550 $Y=1060
X11 8 2 9 11 1 11 8 7 ICV_2 $T=-3665 -3225 0 0 $X=-3120 $Y=1060
X12 9 2 5 3 1 7 3 10 ICV_2 $T=-1235 -3225 0 0 $X=-690 $Y=1060
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4
** N=5 EP=4 IP=8 FDC=60
X0 3 1 4 2 DFF $T=0 0 0 0 $X=-5550 $Y=1060
X1 3 1 4 5 DFF $T=9640 0 0 0 $X=4090 $Y=1060
.ENDS
***************************************
.SUBCKT NAND_0 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT MUX 1 2 3 4
** N=9 EP=4 IP=19 FDC=14
X0 1 3 6 2 INVERTER $T=6025 2225 0 0 $X=7635 $Y=2225
X1 4 1 3 5 7 NAND_0 $T=3445 -2060 0 0 $X=3990 $Y=2225
X2 7 1 3 8 2 NAND_0 $T=4660 -2060 0 0 $X=5205 $Y=2225
X3 5 1 3 9 6 NAND_0 $T=5875 -2060 0 0 $X=6420 $Y=2225
.ENDS
***************************************
.SUBCKT INPUT
** N=11 EP=0 IP=48 FDC=356
X4 10 5 11 1 DFF $T=43985 2105 0 0 $X=38435 $Y=3165
X5 10 5 11 2 DFF $T=58275 2105 0 0 $X=52725 $Y=3165
X6 10 5 11 3 DFF $T=72565 2105 0 0 $X=67015 $Y=3165
X7 10 5 11 6 DFF $T=144695 2105 0 0 $X=139145 $Y=3165
X8 5 4 10 11 ICV_3 $T=86855 2105 0 0 $X=81305 $Y=3165
X9 5 7 10 11 ICV_3 $T=106135 2105 0 0 $X=100585 $Y=3165
X10 5 8 10 11 ICV_3 $T=125415 2105 0 0 $X=119865 $Y=3165
X11 10 9 5 1 MUX $T=42295 940 1 180 $X=33780 $Y=3165
X12 10 9 5 2 MUX $T=56585 940 1 180 $X=48070 $Y=3165
X13 10 9 5 3 MUX $T=70875 940 1 180 $X=62360 $Y=3165
X14 10 9 5 4 MUX $T=85165 940 1 180 $X=76650 $Y=3165
.ENDS
***************************************
