* SPICE NETLIST
***************************************

.SUBCKT M1_N_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_P_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT M1_POLY_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_vtg_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=2
M0 5 1 3 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=2.282e-13 AS=1.834e-13 PD=3.54e-06 PS=3.49e-06 $X=0 $Y=0 $D=5
M1 4 2 5 4 NMOS_VTG L=5e-08 W=1.63e-06 AD=1.77425e-13 AS=2.282e-13 PD=3.485e-06 PS=3.54e-06 $X=380 $Y=0 $D=5
.ENDS
***************************************
.SUBCKT pmos_vtg_0 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 3 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=2.016e-13 AS=1.512e-13 PD=3.16e-06 PS=3.11e-06 $X=0 $Y=0 $D=4
M1 3 2 4 3 PMOS_VTG L=5e-08 W=1.44e-06 AD=1.58175e-13 AS=2.016e-13 PD=3.105e-06 PS=3.16e-06 $X=380 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT NAND 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT MUX 1 2 3 4 5 6
** N=9 EP=6 IP=31 FDC=14
M0 8 2 1 1 NMOS_VTG L=5e-08 W=1.44e-06 AD=1.161e-13 AS=1.0845e-13 PD=3.36e-06 PS=3.19e-06 $X=8070 $Y=2335 $D=5
M1 8 2 3 3 PMOS_VTG L=5e-08 W=1.96e-06 AD=1.6015e-13 AS=1.57e-13 PD=4.57e-06 PS=4.5e-06 $X=8065 $Y=5565 $D=4
X18 4 1 3 7 9 NAND $T=3445 -2060 0 0 $X=3990 $Y=2225
X19 9 1 3 5 2 NAND $T=4660 -2060 0 0 $X=5205 $Y=2225
X20 7 1 3 6 8 NAND $T=5875 -2060 0 0 $X=6420 $Y=2225
.ENDS
***************************************
.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=12 FDC=28
X0 3 9 2 1 4 5 MUX $T=0 0 0 0 $X=3990 $Y=2225
X1 3 10 2 6 7 8 MUX $T=4650 0 0 0 $X=8640 $Y=2225
.ENDS
***************************************
.SUBCKT NAND_0 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=4
X2 4 5 1 2 nmos_vtg_1 $T=945 4395 0 0 $X=695 $Y=4285
X3 4 5 3 1 pmos_vtg_0 $T=945 8045 0 0 $X=695 $Y=7935
.ENDS
***************************************
.SUBCKT MULT
** N=25 EP=0 IP=88 FDC=176
X0 6 17 16 4 5 6 MUX $T=6560 -1025 0 0 $X=10550 $Y=1200
X1 6 17 16 15 6 10 MUX $T=50840 -1025 0 0 $X=54830 $Y=1200
X14 19 16 6 4 1 1 2 3 7 24 ICV_3 $T=-2740 -1025 0 0 $X=1250 $Y=1200
X15 20 16 6 9 8 8 6 5 25 7 ICV_3 $T=12425 -1025 0 0 $X=16415 $Y=1200
X16 9 16 6 2 10 21 12 11 17 25 ICV_3 $T=21725 -1025 0 0 $X=25715 $Y=1200
X17 11 16 6 6 10 12 5 3 13 17 ICV_3 $T=31025 -1025 0 0 $X=35015 $Y=1200
X18 22 16 6 15 14 14 3 2 13 24 ICV_3 $T=41540 -1025 0 0 $X=45530 $Y=1200
X19 7 6 16 17 18 NAND_0 $T=14655 -3085 0 0 $X=15200 $Y=1200
X20 13 6 16 18 23 NAND_0 $T=43770 -3085 0 0 $X=44315 $Y=1200
.ENDS
***************************************
